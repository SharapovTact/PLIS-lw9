----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:24:26 12/15/2025 
-- Design Name: 
-- Module Name:    INVERTOR_7_to_0 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity INVERTOR_7_to_0 is
    Port ( INPUT : in  STD_LOGIC_VECTOR (7 downto 0);
           OUTPUT : in  STD_LOGIC_VECTOR (7 downto 0));
end INVERTOR_7_to_0;

architecture Behavioral of INVERTOR_7_to_0 is

begin
	OUTPUT <= not(INPUT);
	
end Behavioral;

